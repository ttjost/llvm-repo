library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use work.rvex_pkg.all;

entity i_mem is
  generic (
    ISSUE_WIDTH : natural := 4);
  port ( 
    clk         : in std_logic;
    clk_enable  : in std_logic;
    address     : in std_logic_vector(ADDR_WIDTH - 1 downto 0);     -- address of instruction to be read
    instruction : out std_logic_vector(32*ISSUE_WIDTH - 1 downto 0) 	-- instruction (4 syllables)
  );
end entity i_mem;

architecture rtl of i_mem is
  signal instr : std_logic_vector(32*ISSUE_WIDTH - 1 downto 0) := (others => '0');
begin

  instruction <= instr;

  memory : process(clk)
  begin
    if clk'event and clk = '1' and clk_enable = '1' then
      case address is
        when "0000000000000" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000100000100010000000010000000"&
          "10010000000001001000001001100010";
        when "0000000000001" => instr <=
          "10000010000000000000000000100010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000000010" => instr <=
          "00000010000000000000000000101000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000000011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000000100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000011111000001001100010";
        when "0000000000101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000000110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000000111" => instr <=
          "10110010000010001111001000010101"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000001000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000001001" => instr <=
          "10100010000010001111010000010101"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000001010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000001011" => instr <=
          "10010010000010001111011000010101"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000001100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000001101" => instr <=
          "10000010000010001111100000010101"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000001110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000001111" => instr <=
          "01110010000010001111101000010101"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000010000" => instr <=
          "01110000000001001111101001100010"&
          "00101000000000001111100001100010"&
          "00000000000100000000000010000000"&
          "10010000000001001000011001100010";
        when "0000000010001" => instr <=
          "01100010000010001000000000001110"&
          "00000100000100000000000010001010"&
          "01010000000001001111011001100010"&
          "00000100000100000000000010000110";
        when "0000000010010" => instr <=
          "00000000000000000000000001100000"&
          "01100000000001110000110001100010"&
          "10000000000001110000101001100010"&
          "10100000000001110000100001100010";
        when "0000000010011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000010100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000001011100000000000100010";
        when "0000000010101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000010110" => instr <=
          "00000100000100000000000010000100"&
          "00000000000001001111001001100010"&
          "00000100000100000000000010000000"&
          "01100000000001001111010001100010";
        when "0000000010111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10100000000001110000011001100010";
        when "0000000011000" => instr <=
          "00000000000000000000000001100000"&
          "01000000000001110000110001100010"&
          "10000000000001110000101001100010"&
          "00100000000001110000100001100010";
        when "0000000011001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000011010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000010001000000000000100010";
        when "0000000011011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000011100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11110100000001111001011001100010";
        when "0000000011101" => instr <=
          "00000010110110001001100100010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000011110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000011111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000100000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10000000011000001000000001010011";
        when "0000000100001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000100010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000100011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000100100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10000000001001100000000000100100";
        when "0000000100101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000100110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000100111" => instr <=
          "00001010110110001001100100010011"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000101000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000101001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000101010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000011000000001100000011101";
        when "0000000101011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000101100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000100011000001000000001010011";
        when "0000000101101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000101110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000101111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000110000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10000000001000110000000000100100";
        when "0000000110001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000110010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11111000000001111001011001100010";
        when "0000000110011" => instr <=
          "00000010110100001001100100010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000110100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000110101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000110110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10000000011000001000000001010011";
        when "0000000110111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000111000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000111001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000111010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000001000010000000000100100";
        when "0000000111011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000111100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000111101" => instr <=
          "00001010110100001001100100010011"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000111110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000000111111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001000000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000011000000001100000011101";
        when "0000001000001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001000010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000100011000001000000001010011";
        when "0000001000011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001000100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001000101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001000110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000111100000000000100100";
        when "0000001000111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001001000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000001001011001100010"&
          "00000000000100000000000010000000"&
          "00000000000001011001100001100010";
        when "0000001001001" => instr <=
          "00000010110010001001101100010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001001010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001001011" => instr <=
          "00000010011000001001110000010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001001100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001001101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001001110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11000000011010010000000001010011";
        when "0000001001111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001010000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001010001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001010010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000110110000000000100100";
        when "0000001010011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001010100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000100000000001001011001100010";
        when "0000001010101" => instr <=
          "00001010110010001001101100010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001010110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001010111" => instr <=
          "00001010011000001001110000010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001011000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001011001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001011010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11000000011010010000000001000001";
        when "0000001011011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001011100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001011101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001011110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000110000000000000100101";
        when "0000001011111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001100000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00001000000000001001011001100010";
        when "0000001100001" => instr <=
          "00010010110010001001101100010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001100010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001100011" => instr <=
          "00010010011000001001110000010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001100100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001100101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001100110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11000000011010010000000001010011";
        when "0000001100111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001101000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001101001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001101010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000101010000000000100100";
        when "0000001101011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001101100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00001100000000001001011001100010";
        when "0000001101101" => instr <=
          "00011010110010001001101100010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001101110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001101111" => instr <=
          "00011010011000001001110000010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001110000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001110001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001110010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11000000011010010000000001010011";
        when "0000001110011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001110100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001110101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001110110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000100100000000000100100";
        when "0000001110111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001111000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00010000000000001001011001100010";
        when "0000001111001" => instr <=
          "00100010110010001001101100010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001111010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001111011" => instr <=
          "00100010011000001001110000010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001111100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001111101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000001111110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11000000011010010000000001010011";
        when "0000001111111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010000000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010000001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010000010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000011110000000000100100";
        when "0000010000011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010000100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00010100000000001001011001100010";
        when "0000010000101" => instr <=
          "00101010110010001001101100010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010000110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010000111" => instr <=
          "00101010011000001001110000010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010001000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010001001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010001010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11000000011010010000000001010011";
        when "0000010001011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010001100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010001101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010001110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000011000000000000100100";
        when "0000010001111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010010000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00011000000000001001011001100010";
        when "0000010010001" => instr <=
          "00110010110010001001101100010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010010010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010010011" => instr <=
          "00110010011000001001110000010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010010100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010010101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010010110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11000000011010010000000001010011";
        when "0000010010111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010011000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010011001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010011010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000010010000000000100100";
        when "0000010011011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010011100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00011100000000001001011001100010";
        when "0000010011101" => instr <=
          "00111010110010001001101100010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010011110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010011111" => instr <=
          "00111010011000001001110000010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010100000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010100001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010100010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11000000011010010000000001010011";
        when "0000010100011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010100100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010100101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010100110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000001100000000000100100";
        when "0000010100111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010101000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00100000000000001001011001100010";
        when "0000010101001" => instr <=
          "01000010110010001001101100010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010101010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010101011" => instr <=
          "01000010011000001001110000010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010101100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010101101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010101110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11000000011010010000000001010011";
        when "0000010101111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010110000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010110001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010110010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000110000000000100100";
        when "0000010110011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010110100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11111100000001111001011001100010";
        when "0000010110101" => instr <=
          "01001010110010001001101100010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010110110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010110111" => instr <=
          "01001010011000001001100000010010"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010111000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010111001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010111010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10000000011010010000000001000001";
        when "0000010111011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010111100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010111101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000010111110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00100100010110001000011000111000"&
          "10000000000000000000000000100000";
        when "0000010111111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011000000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "01100000000000010000011001100010";
        when "0000011000001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011000010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011000011" => instr <=
          "01100010000010001000000000001101"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011000100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011000101" => instr <=
          "01110010000010001111101000010000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011000110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011000111" => instr <=
          "10000010000010001111100000010000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011001000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011001001" => instr <=
          "10010010000010001111011000010000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011001010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011001011" => instr <=
          "10100010000010001111010000010000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011001100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000001000010000000000000100110";
        when "0000011001101" => instr <=
          "10110010000010001111001000010000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011001110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011001111" => instr <=
          "00001010001100001001011000010011"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011010000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000100001010001000000001001111";
        when "0000011010001" => instr <=
          "00000010001100001001111000010001"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011010010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011010011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011010100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10000000000101000000000000100100";
        when "0000011010101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011010110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000100000000000010000000"&
          "01010000000001011001100001100010";
        when "0000011010111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011011000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10000000010110010001101001101100";
        when "0000011011001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011011010" => instr <=
          "00000000000000001010001001100010"&
          "01111100000000001010000001100010"&
          "00000100000000001001110001100010"&
          "00000100001010001001101001100010";
        when "0000011011011" => instr <=
          "00000010011010001011011000010000"&
          "00000000000000000000000001100000"&
          "00001000000000001010011001100010"&
          "00001100000000001010010001100010";
        when "0000011011100" => instr <=
          "11111100000000000000000010000100"&
          "11111100000001111010101001100010"&
          "00000100000100000000000010000000"&
          "11100000000000101010100001100010";
        when "0000011011101" => instr <=
          "01100010000000000011001001100010"&
          "10000000000000000011000001100010"&
          "11000000000000010011010001100010"&
          "00010000000000001010111001100010";
        when "0000011011110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011011111" => instr <=
          "00000010110010001011100000010001"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011100000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011100001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011100010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10000000011110110011100000011010";
        when "0000011100011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011100100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000111000100011101000011000";
        when "0000011100101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011100110" => instr <=
          "00100000111010001011110001100011"&
          "11000000110110010100001000011000"&
          "01000000110110100100000000011000"&
          "10100000111000110011111001100010";
        when "0000011100111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011101000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10100000111110110100010000011111";
        when "0000011101001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011101010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "01100000000100110000000101001111";
        when "0000011101011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011101100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011101101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011101110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00010000100010001011111000111000"&
          "01100000100010110100011000111000";
        when "0000011101111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011110000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "01000000000111000100000100011010"&
          "00000000000111000011101101100010";
        when "0000011110001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011110010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00100000000001000000000101001111";
        when "0000011110011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011110100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011110101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011110110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10000000000000000000000000100100";
        when "0000011110111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011111000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000011000100000100011010"&
          "00100000111011000011101001100010"&
          "00001000111110001011111001101001";
        when "0000011111001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011111010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "01100000110110100100001000011000";
        when "0000011111011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011111100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11000000111110110011011001101001"&
          "00100000000001000000000101000011";
        when "0000011111101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011111110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000011111111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100000000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00100000000001000000000101001111"&
          "00000100000000001011110000110000";
        when "0000100000001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100000010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11000000110110110011011001101001";
        when "0000100000011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100000100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10000000110110100011111001101100"&
          "00100000100011000011110000111000";
        when "0000100000101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100000110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11111100111001111000000001000111"&
          "10100000111100110011101001100010";
        when "0000100000111" => instr <=
          "00000010111110001011100000010000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100001000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00100000111010100011110000011010";
        when "0000100001001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100001010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11000000111010110011100000111000"&
          "01100000111000010001011001100010";
        when "0000100001011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100001100" => instr <=
          "00000000000000000000000001100000"&
          "00000000110100001000000001000001"&
          "00000000010110001001011001100101"&
          "11100000111000010001111001100010";
        when "0000100001101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100001110" => instr <=
          "00000000011110001001111001100101"&
          "11111100000000000000000010000010"&
          "11111100011111111000001001000111"&
          "01100000010110011001011001100111";
        when "0000100001111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000111111111111111110000111";
        when "0000100010000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10000000010110010011010001101100"&
          "00100000000000010000000000100100";
        when "0000100010001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100010010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11100000110110100010110001101111";
        when "0000100010011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100010100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000101100000010110000011101"&
          "10100000000000010000000000100000";
        when "0000100010101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100010110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00111100110110001011011001100011";
        when "0000100010111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100011000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000100110000001011100001100010"&
          "11000000110110100011011001101001";
        when "0000100011001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100011010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10000000000000110011000001100010";
        when "0000100011011" => instr <=
          "00000010110000001011011000010111"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100011100" => instr <=
          "00000100000000001011010000110000"&
          "11111100011011111001101001100010"&
          "11100000101010010001111000111001"&
          "00001000110010001011001001100010";
        when "0000100011101" => instr <=
          "00000010110100001011011000010000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100011110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000100011010001000001001000111";
        when "0000100011111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100100000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100100001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100100010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10100100111011101111111100100100";
        when "0000100100011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100100100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10100000000000000000000000100100";
        when "0000100100101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100100110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100100111" => instr <=
          "00000010110000001010110000010111"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100101000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100101001" => instr <=
          "00000010001100001001111000010110"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100101010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000001000000000000000000100110";
        when "0000100101011" => instr <=
          "00001010001100001001011000010111"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100101100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100101101" => instr <=
          "00001010001100001001011000010011"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100101110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000100001010001000000001001111";
        when "0000100101111" => instr <=
          "00000010001100001001100000010001"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100110000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100110001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100110010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00100000000011000000000000100100";
        when "0000100110011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100110100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000100000000000010000000"&
          "01010000000001011001101001100010";
        when "0000100110101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100110110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10100000010110010001110001101100";
        when "0000100110111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100111000" => instr <=
          "01111000000000001010001001100010"&
          "01110100000000001010000001100010"&
          "00000000000000001001111001100010"&
          "00000100001010001001110001100010";
        when "0000100111001" => instr <=
          "00000010011100001011001000010000"&
          "01111100000000001010100001100010"&
          "00001100000000001010011001100010"&
          "00000100000000001010010001100010";
        when "0000100111010" => instr <=
          "11111100000001111010111001100010"&
          "00000100000100000000000010000010"&
          "11100000000000101010110001100010"&
          "00001000000000001010101001100010";
        when "0000100111011" => instr <=
          "10000010000000000011100001100010"&
          "11100000000000010011011001100010"&
          "00010000000000001011000001100010"&
          "11111100000000000000000010000110";
        when "0000100111100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "01100000000000000011010001100010";
        when "0000100111101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000100111110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "11000000000000110011101001100010"&
          "00000000110110001000000001010011";
        when "0000100111111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101000000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101000001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101000010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10100000000000010000000000100100";
        when "0000101000011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101000100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000100110100001011010001100010";
        when "0000101000101" => instr <=
          "00000010110100001011101000010011"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101000110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101000111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101001000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000111010110011110000011001";
        when "0000101001001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101001010" => instr <=
          "01100000110010100100010000011000"&
          "01000000110010100100001000011000"&
          "00100000111100100100000001101111"&
          "00000000111100100011111001101111";
        when "0000101001011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00111100111100001100011001100011";
        when "0000101001100" => instr <=
          "11000000000110100100011101101100"&
          "10000000111100100100100001101111"&
          "10000000000000100100000100011000"&
          "10000000111110100011111000011000";
        when "0000101001101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00100000111100001011110001100011"&
          "10100000110010100100101000011000";
        when "0000101001110" => instr <=
          "00000000111100001000000001000001"&
          "00100000000001000100000101100011"&
          "10000000001000100011111100011000"&
          "00100000111110110011001001100011";
        when "0000101001111" => instr <=
          "00000010000110001100001100010000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101010000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10100000111111000011110001100011"&
          "01000000110011000011001001100010";
        when "0000101010001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101010010" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000110011000011001001100010"&
          "01100000000010010001011101100010";
        when "0000101010011" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101010100" => instr <=
          "00000000000000000000000001100000"&
          "11000000110010110011001001100010"&
          "00000000110110001000001001000001"&
          "00000000010110001001011001100101";
        when "0000101010101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101010110" => instr <=
          "00000000000000000000000001100000"&
          "11100000110010010011011000011010"&
          "11111100011101111001110001100010"&
          "01100000010110011001011001100111";
        when "0000101010111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101011000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "01100000110010110011011000111000"&
          "10100000010110010011110001101100";
        when "0000101011001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101011010" => instr <=
          "00000100000000001011011000110001"&
          "00000100011100001000000001000111"&
          "00001000111000001011111001100010"&
          "10000000110110010001100001100010";
        when "0000101011011" => instr <=
          "00000010111100001011001000010000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101011100" => instr <=
          "00000000111111111111111110000101"&
          "00000000011000001001100001100101"&
          "11111100000000000000000010000000"&
          "11111100011001111000001001000111";
        when "0000101011101" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101011110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101011111" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101100000" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "10000000101110010001100000111001";
        when "0000101100001" => instr <=
          "00000010000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101100010" => instr <=
          "00000000000000000000000001100000"&
          "11100000000000110011100001100010"&
          "10100000000000110011110001100010"&
          "10100000111101101111111100100100";
        when "0000101100011" => instr <=
          "00000010111000001001100000010110"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101100100" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101100101" => instr <=
          "00000010001100001001100000010110"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";
        when "0000101100110" => instr <=
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000001000000000000000000100110";
        when "0000101100111" => instr <=
          "00001010001100001001011000010111"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000"&
          "00000000000000000000000001100000";

        when others  => instr <= (others => '0');
      end case;
    end if;
  end process;

end rtl;
