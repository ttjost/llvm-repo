library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library work;
use work.rVEX_pkg.all;

entity d_mem is
  port (
    clk        : in std_logic; -- system clock
    write_en   : in std_logic_vector(3 downto 0);
    address    : in std_logic_vector((DMEM_LOGDEP - 3) downto 0);
    write_data : in std_logic_vector((DMEM_WIDTH - 1) downto 0);
    read_data  : out std_logic_vector((DMEM_WIDTH - 1) downto 0));
end entity d_mem;

architecture behavioural of d_mem is

  type mem_t is array (0 to (DMEM_DEPTH - 1)) of std_logic_vector((DMEM_WIDTH - 1) downto 0);
  signal d_memory : mem_t := (
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"00000000",
		X"10001000",
		X"18001000",
		X"18001800",
		X"20002000",
		X"00827100",
		X"00000038",
		X"00000000",
		X"11000b00",
		X"17001000",
		X"19001800",
		X"20002100",
		X"07000000",
		X"08000000",
		X"09000000",
		X"0a000000",
		X"0b000000",
		X"0c000000",
		X"0d000000",
		X"0e000000",
		X"10000000",
		X"11000000",
		X"13000000",
		X"15000000",
		X"17000000",
		X"19000000",
		X"1c000000",
		X"1f000000",
		X"22000000",
		X"25000000",
		X"29000000",
		X"2d000000",
		X"32000000",
		X"37000000",
		X"3c000000",
		X"42000000",
		X"49000000",
		X"50000000",
		X"58000000",
		X"61000000",
		X"6b000000",
		X"76000000",
		X"82000000",
		X"8f000000",
		X"9d000000",
		X"ad000000",
		X"be000000",
		X"d1000000",
		X"e6000000",
		X"fd000000",
		X"17010000",
		X"33010000",
		X"51010000",
		X"73010000",
		X"98010000",
		X"c1010000",
		X"ee010000",
		X"20020000",
		X"56020000",
		X"92020000",
		X"d4020000",
		X"1c030000",
		X"6c030000",
		X"c3030000",
		X"24040000",
		X"8e040000",
		X"02050000",
		X"83050000",
		X"10060000",
		X"ab060000",
		X"56070000",
		X"12080000",
		X"e0080000",
		X"c3090000",
		X"bd0a0000",
		X"d00b0000",
		X"ff0c0000",
		X"4c0e0000",
		X"ba0f0000",
		X"4c110000",
		X"07130000",
		X"ee140000",
		X"06170000",
		X"54190000",
		X"dc1b0000",
		X"a51e0000",
		X"b6210000",
		X"15250000",
		X"ca280000",
		X"df2c0000",
		X"5b310000",
		X"4b360000",
		X"b93b0000",
		X"b2410000",
		X"44480000",
		X"7e4f0000",
		X"71570000",
		X"2f600000",
		X"ce690000",
		X"62740000",
		X"ff7f0000",
		X"ffffffff",
		X"ffffffff",
		X"ffffffff",
		X"ffffffff",
		X"02000000",
		X"04000000",
		X"06000000",
		X"08000000",
		X"ffffffff",
		X"ffffffff",
		X"ffffffff",
		X"ffffffff",
		X"02000000",
		X"04000000",
		X"06000000",
		X"08000000",
		others => (others => '0'));
  -- flip-flops to store read adresses
  signal read_addr : std_logic_vector((DMEM_LOGDEP - 3) downto 0):= (others => '0'); 

begin
  mem_handler : process(clk)
  begin
    if (rising_edge(clk)) then
	  for index in 0 to 3 loop
	    if write_en(index) = '1' then
          d_memory(conv_integer(address))((index+1)*8 - 1 downto index*8) <= write_data((index+1)*8 - 1 downto index*8);
		end if;
      end loop;
      read_addr <= address;
    end if;
  end process mem_handler;

  -- combinatorial read data
  read_data <= d_memory(conv_integer(read_addr));

end architecture behavioural;
